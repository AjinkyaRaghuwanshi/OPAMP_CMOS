* OTA symbol
* Defining the OTA schematic here ’ Opamp under test ’
*.subckt Opamp-under-test vinn vinp vout VDD VSS
***************************************************************
.include 180nm_bulk.txt
***************************************************************
*Circuit Description

.param lambda = 90n

* OTA parameters ( to be modified )
.param W1 = 2u
.param W2 = 2u
.param W3 = 2u
.param W4 = 2u
.param W5 = 2u
.param W6 = 2u
.param W7 = 2u
.param W8 = 2u
.param W9 = 2u
.param W10 = 2u
.param W11 = 2u
.param W12 = 2u
.param W13 = 2u
.param W14 = 2u
.param W15 = 2u
.param W16 = 2u
.param W17 = 2u
.param W18 = 2u
.param W19 = 2u
.param W20 = 2u
.param L = 180n
* /OTA parameters ( to be modified )
* OTA schematic (Do not change this )
M1 ip2 vinp in0 VSS nmos L=L W=W1 AS={4*lambda*W1} PS={2*W1+8*lambda} AD={4*lambda*W1} PD={2*W1+8*lambda}
M2 ip1 vinn in0 VSS nmos L=L W=W2 AS={4*lambda*W2} PS={2*W2+8*lambda} AD={4*lambda*W2} PD={2*W2+8*lambda}
M3 in2 vinp ip0 VDD pmos L=L W=W3 AS={4*lambda*W3} PS={2*W3+8*lambda} AD={4*lambda*W3} PD={2*W3+8*lambda}
M4 in1 vinn ip0 VDD pmos L=L W=W4 AS={4*lambda*W4} PS={2*W4+8*lambda} AD={4*lambda*W4} PD={2*W4+8*lambda}
M5 in0 vbn VSS VSS nmos L=L W=W5 AS={4*lambda*W5} PS={2*W5+8*lambda} AD={4*lambda*W5} PD={2*W5+8*lambda}
M6 ip0 vbp VDD VDD pmos L=L W=W6 AS={4*lambda*W6} PS={2*W6+8*lambda} AD={4*lambda*W6} PD={2*W6+8*lambda}
M7 ip1 ip3 VDD VDD pmos L=L W=W7 AS={4*lambda*W7} PS={2*W7+8*lambda} AD={4*lambda*W7} PD={2*W7+8*lambda}
M8 ip2 ip3 VDD VDD pmos L=L W=W8 AS={4*lambda*W8} PS={2*W8+8*lambda} AD={4*lambda*W8} PD={2*W8+8*lambda}
M9 ip3 vb1 ip1 ip1 pmos L=L W=W9 AS={4*lambda*W9} PS={2*W9+8*lambda} AD={4*lambda*W9} PD={2*W9+8*lambda}
M10 ip4 vb1 ip2 ip2 pmos L=L W=W10 AS={4*lambda*W10} PS={2*W10+8*lambda} AD={4*lambda*W10} PD={2*W10+8*lambda}
M11 in3 vb3 ip3 VDD pmos L=L W=W11 AS={4*lambda*W11} PS={2*W11+8*lambda} AD={4*lambda*W11} PD={2*W11+8*lambda}
M12 ip3 vb4 in3 VSS nmos L=L W=W12 AS={4*lambda*W12} PS={2*W12+8*lambda} AD={4*lambda*W12} PD={2*W12+8*lambda}
M13 ip4 vb4 in4 VSS nmos L=L W=W13 AS={4*lambda*W13} PS={2*W13+8*lambda} AD={4*lambda*W13} PD={2*W13+8*lambda}
M14 in4 vb3 ip4 VDD pmos L=L W=W14 AS={4*lambda*W14} PS={2*W14+8*lambda} AD={4*lambda*W14} PD={2*W14+8*lambda}
M15 in3 vb2 in1 VSS nmos L=L W=W15 AS={4*lambda*W15} PS={2*W15+8*lambda} AD={4*lambda*W15} PD={2*W15+8*lambda}
M16 in4 vb2 in2 VSS nmos L=L W=W16 AS={4*lambda*W16} PS={2*W16+8*lambda} AD={4*lambda*W16} PD={2*W16+8*lambda}
M17 in1 in3 VSS VSS nmos L=L W=W17 AS={4*lambda*W17} PS={2*W17+8*lambda} AD={4*lambda*W17} PD={2*W17+8*lambda}
M18 in2 in3 VSS VSS nmos L=L W=W18 AS={4*lambda*W18} PS={2*W18+8*lambda} AD={4*lambda*W18} PD={2*W18+8*lambda}
M19 vout ip4 VDD VDD pmos L=L W=W19 AS={4*lambda*W19} PS={2*W19+8*lambda} AD={4*lambda*W19} PD={2*W19+8*lambda}
M20 vout in4 VSS VSS nmos L=L W=W20 AS={4*lambda*W20} PS={2*W20+8*lambda} AD={4*lambda*W20} PD={2*W20+8*lambda}
Cc1 ip4 vout 4p
Cc2 in4 vout 4p
* /OTA schematic (Do not change this )
***************************************************************
* Adding the load capacitance.
CL vout VSS 5p
* Adding the biasing sources
VBP1 vbp VSS dc 1.28
VBN1 vbn VSS dc 0.5999
VDD1 VDD VSS dc 1.8
VSS1 VSS GND dc 0
VB11 vb1 VSS dc 0.5
VB21 vb2 VSS dc 1.4
VB31 vb3 VSS dc 0.1
VB41 vb4 VSS dc 1.6
* Adding the differential sources
Vdn vinn vx dc 0 ac 0
Vdp vinp vx dc 0 ac 0.4
Vcm vx VSS dc 0.9
* Adding the voltage source for input
**Vi Vir VSS dc 0 ac 0
* Adding resistors for closed loop gain (-1)
**R1 Vir vinn 1k
**R2 vinn vout 1k
***************************************************************
* Control Selection
.control
***************************************************************
* Operating point analysis
op
print all

***************************************************************
* AC analysis
ac dec 100 1 100G
plot v(vout)
plot mag((v(vout))/(v(vinp) - v(vinn)))
plot phase((v(vout))/(v(vinp) - v(vinn)))*180/pi
**measure ac
***************************************************************
* Slew Rate analysis


***************************************************************
* Transient analysis


***************************************************************
* Common Mode DC analysis

***************************************************************
.endc
.end
